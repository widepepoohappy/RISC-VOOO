moduele exec_stage #(
    parameter BITWIDTH = 32,
    parameter NRALUOP = 8
) (



);